module Connect4 (
	input logic clk,
	input logic rst,
	input logic [2:0] column,
	input logic load_btn,
	input logic player,
	output logic [1:0] val0,
	output logic [1:0] val1,
	output logic [1:0] val2,
	output logic [1:0] val3,
	output logic [1:0] val4,
	output logic [1:0] val5
);
	logic swp_player, q_player;
	logic [1:0] mux_out;
	logic en_loading, one_sec, t_out, rst_timer, change;
	logic [28:0] timer;
	logic [3:0] secs;
	
	FSM controller (
		.clk(clk),
		.rst(rst),
		.load(load_btn),
		.time_out(t_out),
		.en_loading(en_loading),
		.rst_timer(rst_timer),
		.change_player(change)
	);
	
	Mux2to1 selector (
		.A(2'b01),	// Value for FPGA player
		.B(2'b10),	// Value for Arduino player
		.S(q_player),
		.Y(mux_out)
	);
	
	Inverter swap (
		.A(q_player),
		.en(change),
		.Y(swp_player)
	);
	
	Counter cycles (
		.clk(clk),
		.rst(rst | rst_timer),
		.en_count(1),
		.count(timer)
	);
	
	Counter seconds (
		.clk(clk),
		.rst(rst | rst_timer),
		.en_count(one_sec),
		.count(secs)
	);
	
	Comparator #(.N(4)) check10secs (
		.A(secs),
		.B(4'd10),
		.cmp(t_out)
	);
	
	Comparator #(.N(26)) check1sec (
		.A(timer),
		.B(26'd49_999_999),
		.cmp(one_sec)
	);
	
	Loader loader (
		.clk(clk),
		.rst(rst),
		.column(column),
		.load(en_loading),
		.mux_out(mux_out),
		.val00(val0),
		.val01(val1),
		.val02(val2),
		.val03(val3),
		.val04(val4),
		.val05(val5)
	);
	
	PlayerRegister current (
		.clk(clk),
		.rst(rst),
		.initial_player(player),
		.D(swp_player),
		.Q(q_player)
	);
	
endmodule

	