module Connect4_tb();

endmodule
