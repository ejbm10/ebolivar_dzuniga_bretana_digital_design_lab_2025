module Inverter (
	input logic A,
	output logic Y
);

	assign Y = ~A;
	
endmodule
